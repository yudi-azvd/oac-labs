module Controlador_multiciclo()



endmodule 
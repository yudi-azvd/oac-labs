module SaidaULA (
	input [31:0] iEntrada.
	output [31:0] oSaida
);

assign oSaida = iEntrada;

endmodule 